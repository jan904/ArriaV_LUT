LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY lock_ff IS
    PORT(
        clk : IN STD_LOGIC;
        rst : IN STD_LOGIC;
        start : IN STD_LOGIC;
        signal_in : IN STD_LOGIC;
        lock : OUT STD_LOGIC
    );
END ENTITY lock_ff;

ARCHITECTURE rtl of lock_ff IS
BEGIN
    PROCESS(clk, rst)
    BEGIN
        IF rst = '1' THEN
            lock <= '0';
        ELSIF rising_edge(clk) THEN
            IF signal_in = '1' THEN
                lock <= '1';
            END IF;
        END IF;
    END PROCESS;
END rtl;